always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	chincoka <= papka;
	artemka_loves <= naked_men;
	artemka_loves <= naked_men
	artemka_loves <= naked_men
	artemka_loves <= naked_men
	
end