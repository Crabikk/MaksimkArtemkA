always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
<<<<<<< HEAD
	chincoka <= papka;
=======
	artemka_loves <= naked_men
>>>>>>> 757cdc6fb54c773530b776e07cfce4dd98c2c036
end