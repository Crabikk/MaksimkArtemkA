always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	chincoka <= papka;
	artemka_loves <= naked_men;
	maksimka_loves <= candies;
end