always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	artemka <= loves_naked_men
	chincoka <= papka;
	artemka_loves <= naked_men;
	maksimka_loves <= candies;
end