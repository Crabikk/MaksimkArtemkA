always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	chincoka <= papka;
end