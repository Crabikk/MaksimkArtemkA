always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	artemka_loves <= naked_men
end