always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
<<<<<<< HEAD
	artemka <= loves_naked_men
	chincoka <= papka;
	artemka_loves <= naked_men;
	maksimka_loves <= candies;
=======
	chincoka <= papka;
	artemka_loves <= naked_men;
	artemka_loves <= naked_men
	artemka_loves <= naked_men
	artemka_loves <= naked_men
	
>>>>>>> dev2
end