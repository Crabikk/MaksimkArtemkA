always_ff@(maksimka) begin
	artemka <= happy
end