always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
end