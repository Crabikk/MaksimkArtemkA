always_ff@(maksimka) begin
	artemka <= happy;
	maksimka <= sad;
	artemka <= loves_naked_men
end